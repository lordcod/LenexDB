<?xml version="1.0" encoding="Windows-1251"?>
<LENEX revisiondate="2024-12-02" created="2024-12-30T11:51:45" version="2.0">
 <MEETS>
  <MEET city="���������" name="������� 1 ���� 2025" course="LCM" reservecount="2" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" nation="RUS" hytek.courseorder="L">
   <AGEDATE value="2025-12-31" type="YEAR" />
   <POOL lanemin="1" lanemax="8" />
   <FACILITY city="���������" nation="RUS" />
   <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
   <SESSIONS>
    <SESSION date="2025-02-09" daytime="09:00" name="800" number="1">
     <EVENTS>
      <EVENT eventid="1059" gender="F" number="1" order="1" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1060" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1063" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1064" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1065" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1066" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1067" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1068" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1069" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1108" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1102" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1080" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1084" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1088" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1099" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1097" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1061" gender="M" number="2" order="2" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1070" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1071" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1072" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1073" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1074" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1075" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1076" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1077" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
     </EVENTS>
    </SESSION>
    <SESSION date="2025-02-09" daytime="12:30" name="2 ������" number="2">
     <EVENTS>
      <EVENT eventid="1206" gender="F" number="3" order="19" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1207" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1208" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1209" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1210" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1211" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1212" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1213" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1214" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1222" gender="M" number="4" order="20" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1223" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1224" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1225" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1226" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1227" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1228" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1229" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1230" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1108" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1102" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1080" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1084" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1088" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1099" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1097" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1238" gender="F" number="5" order="21" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1239" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1240" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1241" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1242" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1243" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1244" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1245" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1246" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1254" gender="M" number="6" order="22" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1255" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1256" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1257" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1258" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1259" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1260" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1261" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1262" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1108" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1102" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1080" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1084" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1088" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1099" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1097" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1270" gender="F" number="7" order="23" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1271" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1272" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1273" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1274" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1275" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1276" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1277" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1278" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1286" gender="M" number="8" order="24" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1287" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1288" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1289" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1290" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1291" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1292" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1293" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1294" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1302" gender="F" number="9" order="25" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1303" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1304" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1305" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1306" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1307" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1308" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1309" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1310" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1318" gender="M" number="10" order="26" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1319" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1320" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1321" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1322" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1323" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1324" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1325" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1326" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1334" gender="F" number="11" order="27" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1335" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1336" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1337" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1338" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1339" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1340" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1341" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1342" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1350" gender="M" number="12" order="28" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1351" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1352" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1353" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1354" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1355" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1356" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1357" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1358" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1366" gender="F" number="13" order="29" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1367" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1368" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1369" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1370" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1371" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1372" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1373" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1374" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1382" gender="M" number="14" order="30" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1383" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1384" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1385" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1386" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1387" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1388" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1389" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1390" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1398" gender="F" number="15" order="31" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1399" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1400" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1401" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1402" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1403" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1404" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1405" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1406" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1414" gender="M" number="16" order="32" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1415" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1416" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1417" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1418" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1419" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1420" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1421" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1422" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1430" gender="F" number="17" order="33" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1431" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1432" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1433" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1434" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1435" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1436" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1437" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1438" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
      <EVENT eventid="1446" gender="M" number="18" order="34" round="TIM" preveventid="-1">
       <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
       <AGEGROUPS>
        <AGEGROUP agegroupid="1447" agemax="9" agemin="9" />
        <AGEGROUP agegroupid="1448" agemax="10" agemin="10" />
        <AGEGROUP agegroupid="1449" agemax="11" agemin="11" />
        <AGEGROUP agegroupid="1450" agemax="12" agemin="12" />
        <AGEGROUP agegroupid="1451" agemax="13" agemin="13" />
        <AGEGROUP agegroupid="1452" agemax="14" agemin="14" />
        <AGEGROUP agegroupid="1453" agemax="15" agemin="15" />
        <AGEGROUP agegroupid="1454" agemax="-1" agemin="16" />
       </AGEGROUPS>
       <TIMESTANDARDREFS>
        <TIMESTANDARDREF marker="��" timestandardlistid="1109" />
        <TIMESTANDARDREF marker="���" timestandardlistid="1104" />
        <TIMESTANDARDREF marker="I" timestandardlistid="1081" />
        <TIMESTANDARDREF marker="II" timestandardlistid="1082" />
        <TIMESTANDARDREF marker="III" timestandardlistid="1087" />
        <TIMESTANDARDREF marker="I��" timestandardlistid="1101" />
        <TIMESTANDARDREF marker="II��" timestandardlistid="1096" />
       </TIMESTANDARDREFS>
      </EVENT>
     </EVENTS>
    </SESSION>
   </SESSIONS>
   <CLUBS>
    <CLUB name="������">
     <CONTACT name="������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="�������" birthdate="2011-02-21" gender="M" athleteid="1" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:50.00" />
        <ENTRY eventid="1414" entrytime="03:00:35.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2010-02-16" gender="M" athleteid="2" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:13.22" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="������" birthdate="2013-05-21" gender="M" athleteid="27">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:30.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������������" firstname="������" birthdate="2013-05-22" gender="F" athleteid="36" license="I��">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:000:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="�����" birthdate="2014-03-17" gender="F" athleteid="38">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:13:14.90" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2011-07-03" gender="M" athleteid="48" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:07.26" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="�����" birthdate="2011-02-22" gender="M" athleteid="51" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�����������" firstname="������" birthdate="2012-12-02" gender="M" athleteid="52">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:50.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�� ������">
     <CONTACT name="�� ������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="������" birthdate="2011-08-03" gender="M" athleteid="3" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:45.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="������">
     <CONTACT name="������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2014-08-19" gender="M" athleteid="4" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:14.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�������� �� �����">
     <CONTACT name="�������� �� �����" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2013-03-22" gender="M" athleteid="5" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:25.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�� &quot;�����&quot; �������">
     <CONTACT name="�� &quot;�����&quot; �������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="������" birthdate="2013-08-07" gender="M" athleteid="6" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:09.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���������" firstname="���������" birthdate="2012-10-07" gender="F" athleteid="9" license="II">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:11:05.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="������" birthdate="2013-12-14" gender="M" athleteid="12">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���������" firstname="�����" birthdate="2012-05-17" gender="F" athleteid="13">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:10:23.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="������" birthdate="2009-05-14" gender="M" athleteid="15">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:09:43.95" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="������" birthdate="2012-05-12" gender="M" athleteid="39" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:14.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="������" birthdate="2015-09-24" gender="M" athleteid="40" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�����" firstname="����" birthdate="2012-05-27" gender="M" athleteid="95" license="I">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:09:38.84" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�� ���������� �������">
     <CONTACT name="�� ���������� �������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="������" birthdate="2014-08-14" gender="M" athleteid="7">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:13:16.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������������" firstname="������" birthdate="2011-10-07" gender="F" athleteid="10" license="I��">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:14:04.15" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="������" birthdate="2011-04-09" gender="M" athleteid="11">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:30.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="������" birthdate="2011-04-15" gender="M" athleteid="16" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:37.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���������" firstname="�������" birthdate="2010-08-13" gender="M" athleteid="19">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:55.57" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2012-04-09" gender="F" athleteid="20">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:13:05.41" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="������" birthdate="2013-06-01" gender="M" athleteid="21">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:59.25" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="���������" birthdate="2012-08-04" gender="M" athleteid="22">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:000:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2014-07-05" gender="F" athleteid="23">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:000:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�����" firstname="����" birthdate="2012-01-27" gender="M" athleteid="24" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:28.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="������" birthdate="2013-08-17" gender="F" athleteid="25">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:13:53.62" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2012-03-06" gender="M" athleteid="37" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:21.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�����" firstname="������" birthdate="2011-07-06" gender="M" athleteid="41" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:09:35.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2013-03-22" gender="M" athleteid="42">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:30.30" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="�������" birthdate="1999-03-01" gender="M" athleteid="43">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�����������" firstname="��������" birthdate="2010-12-01" gender="M" athleteid="44" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:09:36.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="�����" birthdate="2012-12-04" gender="F" athleteid="45">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:11:03.71" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="�������" birthdate="2013-12-30" gender="M" athleteid="46" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:46.63" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="�������" birthdate="2014-06-01" gender="F" athleteid="47">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:12:03.23" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="����" birthdate="2012-04-18" gender="M" athleteid="49">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:06.23" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2010-04-25" gender="F" athleteid="50">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:000:00.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="���� �� ��� ������������">
     <CONTACT name="���� �� ��� ������������" />
     <ATHLETES>
      <ATHLETE lastname="������" firstname="����" birthdate="2014-05-31" gender="F" athleteid="8" license="III">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:13:23.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���������" firstname="�����" birthdate="2014-11-25" gender="F" athleteid="99" license="III">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:12:38.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�������">
     <CONTACT name="�������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="������" birthdate="2014-10-08" gender="M" athleteid="14" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:13:40.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="������������">
     <CONTACT name="������������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="�����" birthdate="2013-09-16" gender="M" athleteid="17" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:14:15.02" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="����" birthdate="2012-02-15" gender="M" athleteid="18" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:14:10.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="������� �����">
     <CONTACT name="������� �����" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="������" birthdate="2013-05-15" gender="F" athleteid="26" license="II">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:11:49.91" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="������">
     <CONTACT name="������" />
     <ATHLETES>
      <ATHLETE lastname="������" firstname="���������" birthdate="2012-03-30" gender="M" athleteid="28" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:03.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="������">
     <CONTACT name="������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="���������" birthdate="2012-05-31" gender="M" athleteid="29">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:55.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� ��ػ �� ����������">
     <CONTACT name="��� ��ػ �� ����������" />
     <ATHLETES>
      <ATHLETE lastname="���������" firstname="����" birthdate="2012-04-04" gender="M" athleteid="30" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:30.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� �� ��� ����">
     <CONTACT name="��� �� ��� ����" />
     <ATHLETES>
      <ATHLETE lastname="������" firstname="������" birthdate="2012-04-27" gender="M" athleteid="31">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:12.89" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2011-09-26" gender="M" athleteid="32">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:23.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="������" birthdate="2013-06-04" gender="M" athleteid="60" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:09.67" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���������" firstname="���������" birthdate="2010-07-22" gender="F" athleteid="80">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:10:30.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2014-01-23" gender="F" athleteid="92">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:14:20.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="������" birthdate="2015-07-15" gender="F" athleteid="94" license="III">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:14:10.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="����" birthdate="2013-12-15" gender="M" athleteid="97" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:51.62" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��������">
     <CONTACT name="��������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="�����" birthdate="2014-01-06" gender="M" athleteid="33" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:44.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="Vpride">
     <CONTACT name="Vpride" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="��������" birthdate="2015-04-18" gender="M" athleteid="34">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:40.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="���������">
     <CONTACT name="���������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="������" birthdate="2012-01-05" gender="M" athleteid="35" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:35.80" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���" firstname="��������" birthdate="2010-04-28" gender="M" athleteid="61" license="I">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:08:58.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="���������" birthdate="2012-06-18" gender="M" athleteid="70">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:50.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="����" firstname="������" birthdate="2012-08-21" gender="M" athleteid="71" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:13:17.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�K BOGDANOV_TEAM">
     <CONTACT name="�K BOGDANOV_TEAM" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2014-02-09" gender="M" athleteid="53" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:30.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�� ������������">
     <CONTACT name="�� ������������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="�����" birthdate="2010-12-02" gender="M" athleteid="54" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:30.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="������">
     <CONTACT name="������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2011-05-14" gender="M" athleteid="55">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:09:40.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="����� ����� ������">
     <CONTACT name="����� ����� ������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="������" birthdate="2012-05-28" gender="M" athleteid="56" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:30.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="������������">
     <CONTACT name="������������" />
     <ATHLETES>
      <ATHLETE lastname="����������" firstname="�������" birthdate="2013-01-11" gender="M" athleteid="57">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:13:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="����������" birthdate="2014-10-16" gender="F" athleteid="62" license="I��">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:15:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="����" birthdate="2011-03-31" gender="M" athleteid="82" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:14:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="�����" birthdate="2011-06-16" gender="M" athleteid="84">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:10.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="������" birthdate="2014-08-19" gender="F" athleteid="85" license="I��">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:15:40.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2010-11-08" gender="M" athleteid="86">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:15.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="��������" birthdate="2011-06-15" gender="M" athleteid="87" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:00.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="�������" birthdate="2011-06-15" gender="M" athleteid="88" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:30.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="������" birthdate="2010-02-21" gender="M" athleteid="89">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:30.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="����" birthdate="2011-07-25" gender="M" athleteid="90" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:30.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="����� �� &quot;������������&quot;">
     <CONTACT name="����� �� &quot;������������&quot;" />
     <ATHLETES>
      <ATHLETE lastname="���������" firstname="����" birthdate="2010-11-22" gender="M" athleteid="58" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:50.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�������������">
     <CONTACT name="�������������" />
     <ATHLETES>
      <ATHLETE lastname="����������" firstname="�����" birthdate="2011-10-07" gender="M" athleteid="59" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:35.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���������" firstname="��������" birthdate="2010-08-20" gender="M" athleteid="79" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:35.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��������">
     <CONTACT name="��������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="����" birthdate="2012-04-03" gender="M" athleteid="63" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:55.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2015-04-20" gender="M" athleteid="64" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:05.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="����� �� ������, ���������">
     <CONTACT name="����� �� ������, ���������" />
     <ATHLETES>
      <ATHLETE lastname="����������" firstname="����" birthdate="2013-10-25" gender="M" athleteid="65" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:13:09.60" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="������" firstname="����" birthdate="2012-06-13" gender="M" athleteid="67">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:15.85" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="���������" birthdate="2012-05-19" gender="M" athleteid="74" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:33.31" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�������">
     <CONTACT name="�������" />
     <ATHLETES>
      <ATHLETE lastname="�����������" firstname="���������" birthdate="2011-11-11" gender="M" athleteid="66" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:40.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� �� �� ����� (������� �.�)">
     <CONTACT name="��� �� �� ����� (������� �.�)" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2012-11-20" gender="M" athleteid="68" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:48.90" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="����" birthdate="2013-08-12" gender="M" athleteid="69" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:29.50" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="���������" firstname="��������" birthdate="2012-11-16" gender="F" athleteid="75" license="III">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:12:25.80" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="������" birthdate="2013-07-04" gender="M" athleteid="76" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:59.90" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�����" birthdate="2012-01-29" gender="M" athleteid="77" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:09:55.80" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="������" birthdate="2013-01-23" gender="F" athleteid="78" license="II">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:11:15.30" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� �� &quot;���� �� ��������&quot; ������">
     <CONTACT name="��� �� &quot;���� �� ��������&quot; ������" />
     <ATHLETES>
      <ATHLETE lastname="��������" firstname="���������" birthdate="2013-06-14" gender="M" athleteid="72" license="II">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:10:50.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2012-12-07" gender="M" athleteid="73" license="III">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:07.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2012-07-21" gender="M" athleteid="93">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:18.50" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="�������">
     <CONTACT name="�������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="������" birthdate="2012-03-02" gender="F" athleteid="81" license="I">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:10:10.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="���������">
     <CONTACT name="���������" />
     <ATHLETES>
      <ATHLETE lastname="������" firstname="������" birthdate="2014-03-06" gender="M" athleteid="83">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:36.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="����������" firstname="������" birthdate="2014-07-09" gender="M" athleteid="100">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:11:20.00" />
       </ENTRIES>
      </ATHLETE>
      <ATHLETE lastname="��������" firstname="�����" birthdate="2015-09-28" gender="F" athleteid="101" license="I��">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:13:15.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� ������">
     <CONTACT name="��� ������" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="�������" birthdate="2014-06-18" gender="F" athleteid="91" license="III">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:12:00.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� �� &quot;�� &quot;��������&quot;">
     <CONTACT name="��� �� &quot;�� &quot;��������&quot;" />
     <ATHLETES>
      <ATHLETE lastname="�������" firstname="���������" birthdate="2011-07-01" gender="F" athleteid="96" license="II">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:10:27.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� ������">
     <CONTACT name="��� ������" />
     <ATHLETES>
      <ATHLETE lastname="�����" firstname="������" birthdate="2014-06-26" gender="M" athleteid="98" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:12:36.00" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="���������">
     <CONTACT name="���������" />
     <ATHLETES>
      <ATHLETE lastname="���������" firstname="������" birthdate="2013-03-07" gender="F" athleteid="102" license="II">
       <ENTRIES>
        <ENTRY eventid="1059" entrytime="03:11:09.99" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
    <CLUB name="��� �� �� ������ ������� �����">
     <CONTACT name="��� �� �� ������ ������� �����" />
     <ATHLETES>
      <ATHLETE lastname="�����" firstname="�����" birthdate="2011-11-11" gender="M" athleteid="103" license="I��">
       <ENTRIES>
        <ENTRY eventid="1061" entrytime="03:13:10.50" />
       </ENTRIES>
      </ATHLETE>
     </ATHLETES>
    </CLUB>
   </CLUBS>
  </MEET>
 </MEETS>
 <TIMESTANDARDLISTS>
  <TIMESTANDARDLIST timestandardlistid="1078" code="I" course="SCM" gender="F" name="�������� I ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:09.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:53.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:35.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:38.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:10:11.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:52.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:21.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:37.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:03.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:34.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:34.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:20.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:31.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:27.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:20:04.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:13.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:14.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1079" code="I" course="SCM" gender="M" name="�������� I ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:01.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:36.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:31.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:21.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:24.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:25.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:11.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:02.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:56.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:17.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:19.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:05.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.35">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:24.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:05.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:04.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:05.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1080" code="I" course="LCM" gender="F" name="�������� I ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:11.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:56.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:36.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:42.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:10:23.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:59.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:22.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:42.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:05.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:37.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:37.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:23.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:31.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:32.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:28.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:20:27.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:14.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1081" code="I" course="LCM" gender="M" name="�������� I ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:03.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:39.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:32.40">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:25.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:37.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:31.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:13.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:07.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:58.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:20.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:22.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:08.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:27.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:25.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:29.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:06.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1082" code="II" course="LCM" gender="M" name="�������� II ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:11.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:58.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:35.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:44.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:11:14.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:06.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:21.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:48.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:04.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:39.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:38.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:23.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:32.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:27.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:20:50.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:14.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1083" code="II" course="SCM" gender="F" name="�������� II ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:19.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:14.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:40.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:59.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:11:42.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:34.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:29.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:21.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:11.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:55.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:54.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:36.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:33.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:36.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:22:34.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:21.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:23.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1084" code="II" course="LCM" gender="F" name="�������� II ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:20.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:17.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:40.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:03.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:11:54.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:40.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:31.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:27.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:12.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:58.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:57.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:38.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:34.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:37.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:31.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:22:57.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:22.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1085" code="II" course="SCM" gender="M" name="�������� II ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:10.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:55.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:35.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:38.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:11:02.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:00.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:20.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:43.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:03.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:36.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:36.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:20.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:32.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:20:27.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:12.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:13.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1086" code="III" course="SCM" gender="F" name="�������� III ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:30.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:39.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:44.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:25.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:13:15.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:18.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:41.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:14.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:19.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:18.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:16.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:54.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:36.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:40.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:32.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:25:57.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:31.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:34.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1087" code="III" course="LCM" gender="M" name="�������� III ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:21.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:21.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:39.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:08.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:12:36.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:47.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:29.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:37.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:12.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:00.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:59.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:41.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:33.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:36.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:23:50.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:22.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1088" code="III" course="LCM" gender="F" name="�������� III ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:31.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:42.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:44.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:29.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:13:27.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:24.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:43.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:20.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:20.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:21.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:19.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:57.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:37.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:41.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:33.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:26:20.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:32.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1089" code="III" course="SCM" gender="M" name="�������� III ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="9" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:20.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:18.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:38.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:04.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:12:24.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:41.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:28.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:31.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:10.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:57.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:56.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:38.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:33.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:35.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:23:27.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:21.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:23.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1090" code="III�" course="LCM" gender="M" name="�������� III ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:02:10.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:07.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:05.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:48.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:38.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:35.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:24.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:24.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:04.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:39.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:53.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:27.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:58.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:02.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:55.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:35:52.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:17.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1091" code="III�" course="SCM" gender="M" name="�������� III ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:02:01.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:04.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:05.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:44.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:26.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:29.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:23.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:18.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:03.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:36.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:50.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:24.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:58.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:01.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:55.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:35:30.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:16.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:13.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1092" code="III�" course="LCM" gender="F" name="�������� III ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:02:22.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:36.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:12.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:14.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:21:12.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:57.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:38.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:10:43.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:13.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:04.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:18.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:46.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:04.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:07.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:59.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:38:42.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:29.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1093" code="III�" course="SCM" gender="F" name="�������� III ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:02:21.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:33.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:11.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:10.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:21:00.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:51.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:37.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:10:37.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:12.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:01.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:15.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:43.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:03.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:07.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:59.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:38:20.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:28.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:45.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1094" code="II�" course="SCM" gender="F" name="�������� II ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:02:01.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:51.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:01.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:30.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:30.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:40.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:16.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:26.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:53.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:21.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:35.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:05.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:53.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:57.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:49.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:34:10.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:08.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:05.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1095" code="II�" course="SCM" gender="M" name="�������� II ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:49.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:24.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:55.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:04.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:16:26.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:33.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:03.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:22.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:43.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:56.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:10.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:45.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:48.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:51.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:45.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:31:30.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:56.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:53.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1096" code="II�" course="LCM" gender="M" name="�������� II ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:50.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:27.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:55.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:08.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:16:38.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:39.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:04.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:28.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:44.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:59.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:13.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:47.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:48.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:52.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:45.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:31:52.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:57.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1097" code="II�" course="LCM" gender="F" name="�������� II ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:02:02.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:54.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:02.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:34.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:42.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:46.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:17.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:32.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:54.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:24.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:38.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:08.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:54.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:57.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:50.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:34:32.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:09.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1098" code="I�" course="SCM" gender="F" name="�������� I ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:42.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:16.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:51.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:54.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:16:00.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:29.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:06.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:15.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:33.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:45.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:50.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:25.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:43.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:47.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:39.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:30:05.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:45.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:46.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1099" code="I�" course="LCM" gender="F" name="�������� I ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:43.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:19.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:52.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:58.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:16:12.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:35.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:07.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:21.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:34.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:48.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:53.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:28.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:44.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:47.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:40.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:30:27.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:46.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1100" code="I�" course="SCM" gender="M" name="�������� I ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:30.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:51.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:45.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:29.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:14:26.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:37.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:44.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:26.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:23.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:21.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:24.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:04.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:38.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:41.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:35.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:27:30.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:33.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:34.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1101" code="I�" course="LCM" gender="M" name="�������� I ��. ������" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="8" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:31.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:54.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:45.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:33.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:14:38.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:06:43.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:45.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:32.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:24.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:24.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:27.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:07.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:38.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:42.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:35.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:27:52.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:35.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1102" code="���" course="LCM" gender="F" name="�������� ���" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="10" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:06.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:46.40">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:35.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:33.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:42.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:41.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:17.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:20.50">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:01.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:27.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:28.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:14.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:27.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:44.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:10.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1103" code="���" course="SCM" gender="F" name="�������� ���" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="10" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:05.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:43.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:34.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:29.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:30.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:30.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:16.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:15.50">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:00.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:24.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:25.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:11.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:28.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:18:21.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:08.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:09.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1104" code="���" course="LCM" gender="M" name="�������� ���" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="10" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:59.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:29.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:17.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:58.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:14.50">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:08.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:48.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:54.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:13.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:15.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:00.65">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:25.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:28.15">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:23.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:17:29.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:02.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1105" code="���" course="SCM" gender="M" name="�������� ���" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="10" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:58.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:26.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:14.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:50.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:08.50">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:06.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:43.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:53.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:09.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:11.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:57.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:24.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:27.35">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:23.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:17:06.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:00.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:01.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1106" code="��" course="SCM" gender="F" name="�������� ��" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="12" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:01.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:34.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:32.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:20.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:00.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:20.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:12.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:58.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:56.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:16.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:17.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:03.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:27.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:28.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:25.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:17:12.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:03.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:04.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1107" code="��" course="SCM" gender="M" name="�������� ��" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="12" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:54.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:18.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:28.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:05.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:17.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:56.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:03.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:28.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:50.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:02.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:04.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:50.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:23.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:25.89">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:22.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:15:28.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:57.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:56.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1108" code="��" course="LCM" gender="F" name="�������� ��" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="12" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:01:03.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:37.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:33.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:24.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:09:08.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:26.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:13.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:05:03.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:57.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:19.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:20.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:06.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:28.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:17:35.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:06.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1109" code="��" course="LCM" gender="M" name="�������� ��" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="12" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:55.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:21.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:29.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:09.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:25.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:02.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:04.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:34.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:51.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:05.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:07.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:53.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:24.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:23.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:15:51.00">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:58.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1110" code="����" course="SCM" gender="F" name="�������� ����" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="14" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:57.16">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:21.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.04">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:08.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:23.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:03.32">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:05.05">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:35.03">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:52.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:07.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:05.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:55.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:25.62">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:24.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:16:12.06">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:57.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:59.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1111" code="����" course="SCM" gender="M" name="�������� ����" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="14" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:50.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:05.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:54.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:42.70">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:40.94">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:57.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:06.68">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:46.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:52.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:52.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:43.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:22.52">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:23.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:21.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:14:44.74">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:50.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:52.57">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1112" code="����" course="LCM" gender="F" name="�������� ����" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="14" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:58.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:25.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:30.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:12.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:08:31.12">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:08.04">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:06.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:40.80">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:53.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:08.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:09.77">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:56.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:26.03">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:28.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:24.82">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:16:20.88">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:59.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
  <TIMESTANDARDLIST timestandardlistid="1113" code="����" course="LCM" gender="M" name="�������� ����" type="MINIMUM">
   <AGEGROUP agemax="-1" agemin="14" />
   <TIMESTANDARDS>
    <TIMESTANDARD swimtime="00:00:51.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:02:09.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:27.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:58.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:07:52.60">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:03:47.71">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:59.91">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:04:13.76">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:48.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:56.23">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:57.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:01:46.50">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:23.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:24.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:21.92">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:15:06.19">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
    </TIMESTANDARD>
    <TIMESTANDARD swimtime="00:00:53.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
    </TIMESTANDARD>
   </TIMESTANDARDS>
  </TIMESTANDARDLIST>
 </TIMESTANDARDLISTS>
 <CONSTRUCTOR name="Splash ENTRY EDITOR" version="08.00.1343">
  <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
 </CONSTRUCTOR>
</LENEX>
